module dummy_rom(
	input wire [11:0] read_address,
	output reg [7:0] rom_out
);

always @* begin
	case (read_address)
 12'h0: rom_out <= 8'hF0;
 12'h1: rom_out <= 8'h90;
 12'h2: rom_out <= 8'h90;
 12'h3: rom_out <= 8'h90;
 12'h4: rom_out <= 8'hF0;
 12'h5: rom_out <= 8'h20;
 12'h6: rom_out <= 8'h60;
 12'h7: rom_out <= 8'h20;
 12'h8: rom_out <= 8'h20;
 12'h9: rom_out <= 8'h70;
 12'hA: rom_out <= 8'hF0;
 12'hB: rom_out <= 8'h10;
 12'hC: rom_out <= 8'hF0;
 12'hD: rom_out <= 8'h80;
 12'hE: rom_out <= 8'hF0;
 12'hF: rom_out <= 8'hF0;
 12'h10: rom_out <= 8'h10;
 12'h11: rom_out <= 8'hF0;
 12'h12: rom_out <= 8'h10;
 12'h13: rom_out <= 8'hF0;
 12'h14: rom_out <= 8'h90;
 12'h15: rom_out <= 8'h90;
 12'h16: rom_out <= 8'hF0;
 12'h17: rom_out <= 8'h10;
 12'h18: rom_out <= 8'h10;
 12'h19: rom_out <= 8'hF0;
 12'h1A: rom_out <= 8'h80;
 12'h1B: rom_out <= 8'hF0;
 12'h1C: rom_out <= 8'h10;
 12'h1D: rom_out <= 8'hF0;
 12'h1E: rom_out <= 8'hF0;
 12'h1F: rom_out <= 8'h80;
 12'h20: rom_out <= 8'hF0;
 12'h21: rom_out <= 8'h90;
 12'h22: rom_out <= 8'hF0;
 12'h23: rom_out <= 8'hF0;
 12'h24: rom_out <= 8'h10;
 12'h25: rom_out <= 8'h20;
 12'h26: rom_out <= 8'h40;
 12'h27: rom_out <= 8'h40;
 12'h28: rom_out <= 8'hF0;
 12'h29: rom_out <= 8'h90;
 12'h2A: rom_out <= 8'hF0;
 12'h2B: rom_out <= 8'h90;
 12'h2C: rom_out <= 8'hF0;
 12'h2D: rom_out <= 8'hF0;
 12'h2E: rom_out <= 8'h90;
 12'h2F: rom_out <= 8'hF0;
 12'h30: rom_out <= 8'h10;
 12'h31: rom_out <= 8'hF0;
 12'h32: rom_out <= 8'hF0;
 12'h33: rom_out <= 8'h90;
 12'h34: rom_out <= 8'hF0;
 12'h35: rom_out <= 8'h90;
 12'h36: rom_out <= 8'h90;
 12'h37: rom_out <= 8'hE0;
 12'h38: rom_out <= 8'h90;
 12'h39: rom_out <= 8'hE0;
 12'h3A: rom_out <= 8'h90;
 12'h3B: rom_out <= 8'hE0;
 12'h3C: rom_out <= 8'hF0;
 12'h3D: rom_out <= 8'h80;
 12'h3E: rom_out <= 8'h80;
 12'h3F: rom_out <= 8'h80;
 12'h40: rom_out <= 8'hF0;
 12'h41: rom_out <= 8'hE0;
 12'h42: rom_out <= 8'h90;
 12'h43: rom_out <= 8'h90;
 12'h44: rom_out <= 8'h90;
 12'h45: rom_out <= 8'hE0;
 12'h46: rom_out <= 8'hF0;
 12'h47: rom_out <= 8'h80;
 12'h48: rom_out <= 8'hF0;
 12'h49: rom_out <= 8'h80;
 12'h4A: rom_out <= 8'hF0;
 12'h4B: rom_out <= 8'hF0;
 12'h4C: rom_out <= 8'h80;
 12'h4D: rom_out <= 8'hF0;
 12'h4E: rom_out <= 8'h80;
 12'h4F: rom_out <= 8'h80;
 12'h50: rom_out <= 8'h00;
 12'h51: rom_out <= 8'h00;
 12'h52: rom_out <= 8'h00;
 12'h53: rom_out <= 8'h00;
 12'h54: rom_out <= 8'h00;
 12'h55: rom_out <= 8'h00;
 12'h56: rom_out <= 8'h00;
 12'h57: rom_out <= 8'h00;
 12'h58: rom_out <= 8'h00;
 12'h59: rom_out <= 8'h00;
 12'h5A: rom_out <= 8'h00;
 12'h5B: rom_out <= 8'h00;
 12'h5C: rom_out <= 8'h00;
 12'h5D: rom_out <= 8'h00;
 12'h5E: rom_out <= 8'h00;
 12'h5F: rom_out <= 8'h00;
 12'h60: rom_out <= 8'h00;
 12'h61: rom_out <= 8'h00;
 12'h62: rom_out <= 8'h00;
 12'h63: rom_out <= 8'h00;
 12'h64: rom_out <= 8'h00;
 12'h65: rom_out <= 8'h00;
 12'h66: rom_out <= 8'h00;
 12'h67: rom_out <= 8'h00;
 12'h68: rom_out <= 8'h00;
 12'h69: rom_out <= 8'h00;
 12'h6A: rom_out <= 8'h00;
 12'h6B: rom_out <= 8'h00;
 12'h6C: rom_out <= 8'h00;
 12'h6D: rom_out <= 8'h00;
 12'h6E: rom_out <= 8'h00;
 12'h6F: rom_out <= 8'h00;
 12'h70: rom_out <= 8'h00;
 12'h71: rom_out <= 8'h00;
 12'h72: rom_out <= 8'h00;
 12'h73: rom_out <= 8'h00;
 12'h74: rom_out <= 8'h00;
 12'h75: rom_out <= 8'h00;
 12'h76: rom_out <= 8'h00;
 12'h77: rom_out <= 8'h00;
 12'h78: rom_out <= 8'h00;
 12'h79: rom_out <= 8'h00;
 12'h7A: rom_out <= 8'h00;
 12'h7B: rom_out <= 8'h00;
 12'h7C: rom_out <= 8'h00;
 12'h7D: rom_out <= 8'h00;
 12'h7E: rom_out <= 8'h00;
 12'h7F: rom_out <= 8'h00;
 12'h80: rom_out <= 8'h00;
 12'h81: rom_out <= 8'h00;
 12'h82: rom_out <= 8'h00;
 12'h83: rom_out <= 8'h00;
 12'h84: rom_out <= 8'h00;
 12'h85: rom_out <= 8'h00;
 12'h86: rom_out <= 8'h00;
 12'h87: rom_out <= 8'h00;
 12'h88: rom_out <= 8'h00;
 12'h89: rom_out <= 8'h00;
 12'h8A: rom_out <= 8'h00;
 12'h8B: rom_out <= 8'h00;
 12'h8C: rom_out <= 8'h00;
 12'h8D: rom_out <= 8'h00;
 12'h8E: rom_out <= 8'h00;
 12'h8F: rom_out <= 8'h00;
 12'h90: rom_out <= 8'h00;
 12'h91: rom_out <= 8'h00;
 12'h92: rom_out <= 8'h00;
 12'h93: rom_out <= 8'h00;
 12'h94: rom_out <= 8'h00;
 12'h95: rom_out <= 8'h00;
 12'h96: rom_out <= 8'h00;
 12'h97: rom_out <= 8'h00;
 12'h98: rom_out <= 8'h00;
 12'h99: rom_out <= 8'h00;
 12'h9A: rom_out <= 8'h00;
 12'h9B: rom_out <= 8'h00;
 12'h9C: rom_out <= 8'h00;
 12'h9D: rom_out <= 8'h00;
 12'h9E: rom_out <= 8'h00;
 12'h9F: rom_out <= 8'h00;
 12'hA0: rom_out <= 8'h00;
 12'hA1: rom_out <= 8'h00;
 12'hA2: rom_out <= 8'h00;
 12'hA3: rom_out <= 8'h00;
 12'hA4: rom_out <= 8'h00;
 12'hA5: rom_out <= 8'h00;
 12'hA6: rom_out <= 8'h00;
 12'hA7: rom_out <= 8'h00;
 12'hA8: rom_out <= 8'h00;
 12'hA9: rom_out <= 8'h00;
 12'hAA: rom_out <= 8'h00;
 12'hAB: rom_out <= 8'h00;
 12'hAC: rom_out <= 8'h00;
 12'hAD: rom_out <= 8'h00;
 12'hAE: rom_out <= 8'h00;
 12'hAF: rom_out <= 8'h00;
 12'hB0: rom_out <= 8'h00;
 12'hB1: rom_out <= 8'h00;
 12'hB2: rom_out <= 8'h00;
 12'hB3: rom_out <= 8'h00;
 12'hB4: rom_out <= 8'h00;
 12'hB5: rom_out <= 8'h00;
 12'hB6: rom_out <= 8'h00;
 12'hB7: rom_out <= 8'h00;
 12'hB8: rom_out <= 8'h00;
 12'hB9: rom_out <= 8'h00;
 12'hBA: rom_out <= 8'h00;
 12'hBB: rom_out <= 8'h00;
 12'hBC: rom_out <= 8'h00;
 12'hBD: rom_out <= 8'h00;
 12'hBE: rom_out <= 8'h00;
 12'hBF: rom_out <= 8'h00;
 12'hC0: rom_out <= 8'h00;
 12'hC1: rom_out <= 8'h00;
 12'hC2: rom_out <= 8'h00;
 12'hC3: rom_out <= 8'h00;
 12'hC4: rom_out <= 8'h00;
 12'hC5: rom_out <= 8'h00;
 12'hC6: rom_out <= 8'h00;
 12'hC7: rom_out <= 8'h00;
 12'hC8: rom_out <= 8'h00;
 12'hC9: rom_out <= 8'h00;
 12'hCA: rom_out <= 8'h00;
 12'hCB: rom_out <= 8'h00;
 12'hCC: rom_out <= 8'h00;
 12'hCD: rom_out <= 8'h00;
 12'hCE: rom_out <= 8'h00;
 12'hCF: rom_out <= 8'h00;
 12'hD0: rom_out <= 8'h00;
 12'hD1: rom_out <= 8'h00;
 12'hD2: rom_out <= 8'h00;
 12'hD3: rom_out <= 8'h00;
 12'hD4: rom_out <= 8'h00;
 12'hD5: rom_out <= 8'h00;
 12'hD6: rom_out <= 8'h00;
 12'hD7: rom_out <= 8'h00;
 12'hD8: rom_out <= 8'h00;
 12'hD9: rom_out <= 8'h00;
 12'hDA: rom_out <= 8'h00;
 12'hDB: rom_out <= 8'h00;
 12'hDC: rom_out <= 8'h00;
 12'hDD: rom_out <= 8'h00;
 12'hDE: rom_out <= 8'h00;
 12'hDF: rom_out <= 8'h00;
 12'hE0: rom_out <= 8'h00;
 12'hE1: rom_out <= 8'h00;
 12'hE2: rom_out <= 8'h00;
 12'hE3: rom_out <= 8'h00;
 12'hE4: rom_out <= 8'h00;
 12'hE5: rom_out <= 8'h00;
 12'hE6: rom_out <= 8'h00;
 12'hE7: rom_out <= 8'h00;
 12'hE8: rom_out <= 8'h00;
 12'hE9: rom_out <= 8'h00;
 12'hEA: rom_out <= 8'h00;
 12'hEB: rom_out <= 8'h00;
 12'hEC: rom_out <= 8'h00;
 12'hED: rom_out <= 8'h00;
 12'hEE: rom_out <= 8'h00;
 12'hEF: rom_out <= 8'h00;
 12'hF0: rom_out <= 8'h00;
 12'hF1: rom_out <= 8'h00;
 12'hF2: rom_out <= 8'h00;
 12'hF3: rom_out <= 8'h00;
 12'hF4: rom_out <= 8'h00;
 12'hF5: rom_out <= 8'h00;
 12'hF6: rom_out <= 8'h00;
 12'hF7: rom_out <= 8'h00;
 12'hF8: rom_out <= 8'h00;
 12'hF9: rom_out <= 8'h00;
 12'hFA: rom_out <= 8'h00;
 12'hFB: rom_out <= 8'h00;
 12'hFC: rom_out <= 8'h00;
 12'hFD: rom_out <= 8'h00;
 12'hFE: rom_out <= 8'h00;
 12'hFF: rom_out <= 8'h00;
 12'h100: rom_out <= 8'h00;
 12'h101: rom_out <= 8'h00;
 12'h102: rom_out <= 8'h00;
 12'h103: rom_out <= 8'h00;
 12'h104: rom_out <= 8'h00;
 12'h105: rom_out <= 8'h00;
 12'h106: rom_out <= 8'h00;
 12'h107: rom_out <= 8'h00;
 12'h108: rom_out <= 8'h00;
 12'h109: rom_out <= 8'h00;
 12'h10A: rom_out <= 8'h00;
 12'h10B: rom_out <= 8'h00;
 12'h10C: rom_out <= 8'h00;
 12'h10D: rom_out <= 8'h00;
 12'h10E: rom_out <= 8'h00;
 12'h10F: rom_out <= 8'h00;
 12'h110: rom_out <= 8'h00;
 12'h111: rom_out <= 8'h00;
 12'h112: rom_out <= 8'h00;
 12'h113: rom_out <= 8'h00;
 12'h114: rom_out <= 8'h00;
 12'h115: rom_out <= 8'h00;
 12'h116: rom_out <= 8'h00;
 12'h117: rom_out <= 8'h00;
 12'h118: rom_out <= 8'h00;
 12'h119: rom_out <= 8'h00;
 12'h11A: rom_out <= 8'h00;
 12'h11B: rom_out <= 8'h00;
 12'h11C: rom_out <= 8'h00;
 12'h11D: rom_out <= 8'h00;
 12'h11E: rom_out <= 8'h00;
 12'h11F: rom_out <= 8'h00;
 12'h120: rom_out <= 8'h00;
 12'h121: rom_out <= 8'h00;
 12'h122: rom_out <= 8'h00;
 12'h123: rom_out <= 8'h00;
 12'h124: rom_out <= 8'h00;
 12'h125: rom_out <= 8'h00;
 12'h126: rom_out <= 8'h00;
 12'h127: rom_out <= 8'h00;
 12'h128: rom_out <= 8'h00;
 12'h129: rom_out <= 8'h00;
 12'h12A: rom_out <= 8'h00;
 12'h12B: rom_out <= 8'h00;
 12'h12C: rom_out <= 8'h00;
 12'h12D: rom_out <= 8'h00;
 12'h12E: rom_out <= 8'h00;
 12'h12F: rom_out <= 8'h00;
 12'h130: rom_out <= 8'h00;
 12'h131: rom_out <= 8'h00;
 12'h132: rom_out <= 8'h00;
 12'h133: rom_out <= 8'h00;
 12'h134: rom_out <= 8'h00;
 12'h135: rom_out <= 8'h00;
 12'h136: rom_out <= 8'h00;
 12'h137: rom_out <= 8'h00;
 12'h138: rom_out <= 8'h00;
 12'h139: rom_out <= 8'h00;
 12'h13A: rom_out <= 8'h00;
 12'h13B: rom_out <= 8'h00;
 12'h13C: rom_out <= 8'h00;
 12'h13D: rom_out <= 8'h00;
 12'h13E: rom_out <= 8'h00;
 12'h13F: rom_out <= 8'h00;
 12'h140: rom_out <= 8'h00;
 12'h141: rom_out <= 8'h00;
 12'h142: rom_out <= 8'h00;
 12'h143: rom_out <= 8'h00;
 12'h144: rom_out <= 8'h00;
 12'h145: rom_out <= 8'h00;
 12'h146: rom_out <= 8'h00;
 12'h147: rom_out <= 8'h00;
 12'h148: rom_out <= 8'h00;
 12'h149: rom_out <= 8'h00;
 12'h14A: rom_out <= 8'h00;
 12'h14B: rom_out <= 8'h00;
 12'h14C: rom_out <= 8'h00;
 12'h14D: rom_out <= 8'h00;
 12'h14E: rom_out <= 8'h00;
 12'h14F: rom_out <= 8'h00;
 12'h150: rom_out <= 8'h00;
 12'h151: rom_out <= 8'h00;
 12'h152: rom_out <= 8'h00;
 12'h153: rom_out <= 8'h00;
 12'h154: rom_out <= 8'h00;
 12'h155: rom_out <= 8'h00;
 12'h156: rom_out <= 8'h00;
 12'h157: rom_out <= 8'h00;
 12'h158: rom_out <= 8'h00;
 12'h159: rom_out <= 8'h00;
 12'h15A: rom_out <= 8'h00;
 12'h15B: rom_out <= 8'h00;
 12'h15C: rom_out <= 8'h00;
 12'h15D: rom_out <= 8'h00;
 12'h15E: rom_out <= 8'h00;
 12'h15F: rom_out <= 8'h00;
 12'h160: rom_out <= 8'h00;
 12'h161: rom_out <= 8'h00;
 12'h162: rom_out <= 8'h00;
 12'h163: rom_out <= 8'h00;
 12'h164: rom_out <= 8'h00;
 12'h165: rom_out <= 8'h00;
 12'h166: rom_out <= 8'h00;
 12'h167: rom_out <= 8'h00;
 12'h168: rom_out <= 8'h00;
 12'h169: rom_out <= 8'h00;
 12'h16A: rom_out <= 8'h00;
 12'h16B: rom_out <= 8'h00;
 12'h16C: rom_out <= 8'h00;
 12'h16D: rom_out <= 8'h00;
 12'h16E: rom_out <= 8'h00;
 12'h16F: rom_out <= 8'h00;
 12'h170: rom_out <= 8'h00;
 12'h171: rom_out <= 8'h00;
 12'h172: rom_out <= 8'h00;
 12'h173: rom_out <= 8'h00;
 12'h174: rom_out <= 8'h00;
 12'h175: rom_out <= 8'h00;
 12'h176: rom_out <= 8'h00;
 12'h177: rom_out <= 8'h00;
 12'h178: rom_out <= 8'h00;
 12'h179: rom_out <= 8'h00;
 12'h17A: rom_out <= 8'h00;
 12'h17B: rom_out <= 8'h00;
 12'h17C: rom_out <= 8'h00;
 12'h17D: rom_out <= 8'h00;
 12'h17E: rom_out <= 8'h00;
 12'h17F: rom_out <= 8'h00;
 12'h180: rom_out <= 8'h00;
 12'h181: rom_out <= 8'h00;
 12'h182: rom_out <= 8'h00;
 12'h183: rom_out <= 8'h00;
 12'h184: rom_out <= 8'h00;
 12'h185: rom_out <= 8'h00;
 12'h186: rom_out <= 8'h00;
 12'h187: rom_out <= 8'h00;
 12'h188: rom_out <= 8'h00;
 12'h189: rom_out <= 8'h00;
 12'h18A: rom_out <= 8'h00;
 12'h18B: rom_out <= 8'h00;
 12'h18C: rom_out <= 8'h00;
 12'h18D: rom_out <= 8'h00;
 12'h18E: rom_out <= 8'h00;
 12'h18F: rom_out <= 8'h00;
 12'h190: rom_out <= 8'h00;
 12'h191: rom_out <= 8'h00;
 12'h192: rom_out <= 8'h00;
 12'h193: rom_out <= 8'h00;
 12'h194: rom_out <= 8'h00;
 12'h195: rom_out <= 8'h00;
 12'h196: rom_out <= 8'h00;
 12'h197: rom_out <= 8'h00;
 12'h198: rom_out <= 8'h00;
 12'h199: rom_out <= 8'h00;
 12'h19A: rom_out <= 8'h00;
 12'h19B: rom_out <= 8'h00;
 12'h19C: rom_out <= 8'h00;
 12'h19D: rom_out <= 8'h00;
 12'h19E: rom_out <= 8'h00;
 12'h19F: rom_out <= 8'h00;
 12'h1A0: rom_out <= 8'h00;
 12'h1A1: rom_out <= 8'h00;
 12'h1A2: rom_out <= 8'h00;
 12'h1A3: rom_out <= 8'h00;
 12'h1A4: rom_out <= 8'h00;
 12'h1A5: rom_out <= 8'h00;
 12'h1A6: rom_out <= 8'h00;
 12'h1A7: rom_out <= 8'h00;
 12'h1A8: rom_out <= 8'h00;
 12'h1A9: rom_out <= 8'h00;
 12'h1AA: rom_out <= 8'h00;
 12'h1AB: rom_out <= 8'h00;
 12'h1AC: rom_out <= 8'h00;
 12'h1AD: rom_out <= 8'h00;
 12'h1AE: rom_out <= 8'h00;
 12'h1AF: rom_out <= 8'h00;
 12'h1B0: rom_out <= 8'h00;
 12'h1B1: rom_out <= 8'h00;
 12'h1B2: rom_out <= 8'h00;
 12'h1B3: rom_out <= 8'h00;
 12'h1B4: rom_out <= 8'h00;
 12'h1B5: rom_out <= 8'h00;
 12'h1B6: rom_out <= 8'h00;
 12'h1B7: rom_out <= 8'h00;
 12'h1B8: rom_out <= 8'h00;
 12'h1B9: rom_out <= 8'h00;
 12'h1BA: rom_out <= 8'h00;
 12'h1BB: rom_out <= 8'h00;
 12'h1BC: rom_out <= 8'h00;
 12'h1BD: rom_out <= 8'h00;
 12'h1BE: rom_out <= 8'h00;
 12'h1BF: rom_out <= 8'h00;
 12'h1C0: rom_out <= 8'h00;
 12'h1C1: rom_out <= 8'h00;
 12'h1C2: rom_out <= 8'h00;
 12'h1C3: rom_out <= 8'h00;
 12'h1C4: rom_out <= 8'h00;
 12'h1C5: rom_out <= 8'h00;
 12'h1C6: rom_out <= 8'h00;
 12'h1C7: rom_out <= 8'h00;
 12'h1C8: rom_out <= 8'h00;
 12'h1C9: rom_out <= 8'h00;
 12'h1CA: rom_out <= 8'h00;
 12'h1CB: rom_out <= 8'h00;
 12'h1CC: rom_out <= 8'h00;
 12'h1CD: rom_out <= 8'h00;
 12'h1CE: rom_out <= 8'h00;
 12'h1CF: rom_out <= 8'h00;
 12'h1D0: rom_out <= 8'h00;
 12'h1D1: rom_out <= 8'h00;
 12'h1D2: rom_out <= 8'h00;
 12'h1D3: rom_out <= 8'h00;
 12'h1D4: rom_out <= 8'h00;
 12'h1D5: rom_out <= 8'h00;
 12'h1D6: rom_out <= 8'h00;
 12'h1D7: rom_out <= 8'h00;
 12'h1D8: rom_out <= 8'h00;
 12'h1D9: rom_out <= 8'h00;
 12'h1DA: rom_out <= 8'h00;
 12'h1DB: rom_out <= 8'h00;
 12'h1DC: rom_out <= 8'h00;
 12'h1DD: rom_out <= 8'h00;
 12'h1DE: rom_out <= 8'h00;
 12'h1DF: rom_out <= 8'h00;
 12'h1E0: rom_out <= 8'h00;
 12'h1E1: rom_out <= 8'h00;
 12'h1E2: rom_out <= 8'h00;
 12'h1E3: rom_out <= 8'h00;
 12'h1E4: rom_out <= 8'h00;
 12'h1E5: rom_out <= 8'h00;
 12'h1E6: rom_out <= 8'h00;
 12'h1E7: rom_out <= 8'h00;
 12'h1E8: rom_out <= 8'h00;
 12'h1E9: rom_out <= 8'h00;
 12'h1EA: rom_out <= 8'h00;
 12'h1EB: rom_out <= 8'h00;
 12'h1EC: rom_out <= 8'h00;
 12'h1ED: rom_out <= 8'h00;
 12'h1EE: rom_out <= 8'h00;
 12'h1EF: rom_out <= 8'h00;
 12'h1F0: rom_out <= 8'h00;
 12'h1F1: rom_out <= 8'h00;
 12'h1F2: rom_out <= 8'h00;
 12'h1F3: rom_out <= 8'h00;
 12'h1F4: rom_out <= 8'h00;
 12'h1F5: rom_out <= 8'h00;
 12'h1F6: rom_out <= 8'h00;
 12'h1F7: rom_out <= 8'h00;
 12'h1F8: rom_out <= 8'h00;
 12'h1F9: rom_out <= 8'h00;
 12'h1FA: rom_out <= 8'h00;
 12'h1FB: rom_out <= 8'h00;
 12'h1FC: rom_out <= 8'h00;
 12'h1FD: rom_out <= 8'h00;
 12'h1FE: rom_out <= 8'h00;
 12'h1FF: rom_out <= 8'h00;
 12'h200: rom_out <= 8'h00;
 12'h201: rom_out <= 8'hE0;
 12'h202: rom_out <= 8'hA2;
 12'h203: rom_out <= 8'h2A;
 12'h204: rom_out <= 8'h60;
 12'h205: rom_out <= 8'h0C;
 12'h206: rom_out <= 8'h61;
 12'h207: rom_out <= 8'h08;
 12'h208: rom_out <= 8'hD0;
 12'h209: rom_out <= 8'h1F;
 12'h20A: rom_out <= 8'h70;
 12'h20B: rom_out <= 8'h09;
 12'h20C: rom_out <= 8'hA2;
 12'h20D: rom_out <= 8'h39;
 12'h20E: rom_out <= 8'hD0;
 12'h20F: rom_out <= 8'h1F;
 12'h210: rom_out <= 8'hA2;
 12'h211: rom_out <= 8'h48;
 12'h212: rom_out <= 8'h70;
 12'h213: rom_out <= 8'h08;
 12'h214: rom_out <= 8'hD0;
 12'h215: rom_out <= 8'h1F;
 12'h216: rom_out <= 8'h70;
 12'h217: rom_out <= 8'h04;
 12'h218: rom_out <= 8'hA2;
 12'h219: rom_out <= 8'h57;
 12'h21A: rom_out <= 8'hD0;
 12'h21B: rom_out <= 8'h1F;
 12'h21C: rom_out <= 8'h70;
 12'h21D: rom_out <= 8'h08;
 12'h21E: rom_out <= 8'hA2;
 12'h21F: rom_out <= 8'h66;
 12'h220: rom_out <= 8'hD0;
 12'h221: rom_out <= 8'h1F;
 12'h222: rom_out <= 8'h70;
 12'h223: rom_out <= 8'h08;
 12'h224: rom_out <= 8'hA2;
 12'h225: rom_out <= 8'h75;
 12'h226: rom_out <= 8'hD0;
 12'h227: rom_out <= 8'h1F;
 12'h228: rom_out <= 8'h12;
 12'h229: rom_out <= 8'h28;
 12'h22A: rom_out <= 8'hFF;
 12'h22B: rom_out <= 8'h00;
 12'h22C: rom_out <= 8'hFF;
 12'h22D: rom_out <= 8'h00;
 12'h22E: rom_out <= 8'h3C;
 12'h22F: rom_out <= 8'h00;
 12'h230: rom_out <= 8'h3C;
 12'h231: rom_out <= 8'h00;
 12'h232: rom_out <= 8'h3C;
 12'h233: rom_out <= 8'h00;
 12'h234: rom_out <= 8'h3C;
 12'h235: rom_out <= 8'h00;
 12'h236: rom_out <= 8'hFF;
 12'h237: rom_out <= 8'h00;
 12'h238: rom_out <= 8'hFF;
 12'h239: rom_out <= 8'hFF;
 12'h23A: rom_out <= 8'h00;
 12'h23B: rom_out <= 8'hFF;
 12'h23C: rom_out <= 8'h00;
 12'h23D: rom_out <= 8'h38;
 12'h23E: rom_out <= 8'h00;
 12'h23F: rom_out <= 8'h3F;
 12'h240: rom_out <= 8'h00;
 12'h241: rom_out <= 8'h3F;
 12'h242: rom_out <= 8'h00;
 12'h243: rom_out <= 8'h38;
 12'h244: rom_out <= 8'h00;
 12'h245: rom_out <= 8'hFF;
 12'h246: rom_out <= 8'h00;
 12'h247: rom_out <= 8'hFF;
 12'h248: rom_out <= 8'h80;
 12'h249: rom_out <= 8'h00;
 12'h24A: rom_out <= 8'hE0;
 12'h24B: rom_out <= 8'h00;
 12'h24C: rom_out <= 8'hE0;
 12'h24D: rom_out <= 8'h00;
 12'h24E: rom_out <= 8'h80;
 12'h24F: rom_out <= 8'h00;
 12'h250: rom_out <= 8'h80;
 12'h251: rom_out <= 8'h00;
 12'h252: rom_out <= 8'hE0;
 12'h253: rom_out <= 8'h00;
 12'h254: rom_out <= 8'hE0;
 12'h255: rom_out <= 8'h00;
 12'h256: rom_out <= 8'h80;
 12'h257: rom_out <= 8'hF8;
 12'h258: rom_out <= 8'h00;
 12'h259: rom_out <= 8'hFC;
 12'h25A: rom_out <= 8'h00;
 12'h25B: rom_out <= 8'h3E;
 12'h25C: rom_out <= 8'h00;
 12'h25D: rom_out <= 8'h3F;
 12'h25E: rom_out <= 8'h00;
 12'h25F: rom_out <= 8'h3B;
 12'h260: rom_out <= 8'h00;
 12'h261: rom_out <= 8'h39;
 12'h262: rom_out <= 8'h00;
 12'h263: rom_out <= 8'hF8;
 12'h264: rom_out <= 8'h00;
 12'h265: rom_out <= 8'hF8;
 12'h266: rom_out <= 8'h03;
 12'h267: rom_out <= 8'h00;
 12'h268: rom_out <= 8'h07;
 12'h269: rom_out <= 8'h00;
 12'h26A: rom_out <= 8'h0F;
 12'h26B: rom_out <= 8'h00;
 12'h26C: rom_out <= 8'hBF;
 12'h26D: rom_out <= 8'h00;
 12'h26E: rom_out <= 8'hFB;
 12'h26F: rom_out <= 8'h00;
 12'h270: rom_out <= 8'hF3;
 12'h271: rom_out <= 8'h00;
 12'h272: rom_out <= 8'hE3;
 12'h273: rom_out <= 8'h00;
 12'h274: rom_out <= 8'h43;
 12'h275: rom_out <= 8'hE0;
 12'h276: rom_out <= 8'h00;
 12'h277: rom_out <= 8'hE0;
 12'h278: rom_out <= 8'h00;
 12'h279: rom_out <= 8'h80;
 12'h27A: rom_out <= 8'h00;
 12'h27B: rom_out <= 8'h80;
 12'h27C: rom_out <= 8'h00;
 12'h27D: rom_out <= 8'h80;
 12'h27E: rom_out <= 8'h00;
 12'h27F: rom_out <= 8'h80;
 12'h280: rom_out <= 8'h00;
 12'h281: rom_out <= 8'hE0;
 12'h282: rom_out <= 8'h00;
 12'h283: rom_out <= 8'hE0;
 12'h284: rom_out <= 8'h00;
 12'h285: rom_out <= 8'h00;
 12'h286: rom_out <= 8'h00;
 12'h287: rom_out <= 8'h00;
 12'h288: rom_out <= 8'h00;
 12'h289: rom_out <= 8'h00;
 12'h28A: rom_out <= 8'h00;
 12'h28B: rom_out <= 8'h00;
 12'h28C: rom_out <= 8'h00;
 12'h28D: rom_out <= 8'h00;
 12'h28E: rom_out <= 8'h00;
 12'h28F: rom_out <= 8'h00;
 12'h290: rom_out <= 8'h00;
 12'h291: rom_out <= 8'h00;
 12'h292: rom_out <= 8'h00;
 12'h293: rom_out <= 8'h00;
 12'h294: rom_out <= 8'h00;
 12'h295: rom_out <= 8'h00;
 12'h296: rom_out <= 8'h00;
 12'h297: rom_out <= 8'h00;
 12'h298: rom_out <= 8'h00;
 12'h299: rom_out <= 8'h00;
 12'h29A: rom_out <= 8'h00;
 12'h29B: rom_out <= 8'h00;
 12'h29C: rom_out <= 8'h00;
 12'h29D: rom_out <= 8'h00;
 12'h29E: rom_out <= 8'h00;
 12'h29F: rom_out <= 8'h00;
 12'h2A0: rom_out <= 8'h00;
 12'h2A1: rom_out <= 8'h00;
 12'h2A2: rom_out <= 8'h00;
 12'h2A3: rom_out <= 8'h00;
 12'h2A4: rom_out <= 8'h00;
 12'h2A5: rom_out <= 8'h00;
 12'h2A6: rom_out <= 8'h00;
 12'h2A7: rom_out <= 8'h00;
 12'h2A8: rom_out <= 8'h00;
 12'h2A9: rom_out <= 8'h00;
 12'h2AA: rom_out <= 8'h00;
 12'h2AB: rom_out <= 8'h00;
 12'h2AC: rom_out <= 8'h00;
 12'h2AD: rom_out <= 8'h00;
 12'h2AE: rom_out <= 8'h00;
 12'h2AF: rom_out <= 8'h00;
 12'h2B0: rom_out <= 8'h00;
 12'h2B1: rom_out <= 8'h00;
 12'h2B2: rom_out <= 8'h00;
 12'h2B3: rom_out <= 8'h00;
 12'h2B4: rom_out <= 8'h00;
 12'h2B5: rom_out <= 8'h00;
 12'h2B6: rom_out <= 8'h00;
 12'h2B7: rom_out <= 8'h00;
 12'h2B8: rom_out <= 8'h00;
 12'h2B9: rom_out <= 8'h00;
 12'h2BA: rom_out <= 8'h00;
 12'h2BB: rom_out <= 8'h00;
 12'h2BC: rom_out <= 8'h00;
 12'h2BD: rom_out <= 8'h00;
 12'h2BE: rom_out <= 8'h00;
 12'h2BF: rom_out <= 8'h00;
 12'h2C0: rom_out <= 8'h00;
 12'h2C1: rom_out <= 8'h00;
 12'h2C2: rom_out <= 8'h00;
 12'h2C3: rom_out <= 8'h00;
 12'h2C4: rom_out <= 8'h00;
 12'h2C5: rom_out <= 8'h00;
 12'h2C6: rom_out <= 8'h00;
 12'h2C7: rom_out <= 8'h00;
 12'h2C8: rom_out <= 8'h00;
 12'h2C9: rom_out <= 8'h00;
 12'h2CA: rom_out <= 8'h00;
 12'h2CB: rom_out <= 8'h00;
 12'h2CC: rom_out <= 8'h00;
 12'h2CD: rom_out <= 8'h00;
 12'h2CE: rom_out <= 8'h00;
 12'h2CF: rom_out <= 8'h00;
 12'h2D0: rom_out <= 8'h00;
 12'h2D1: rom_out <= 8'h00;
 12'h2D2: rom_out <= 8'h00;
 12'h2D3: rom_out <= 8'h00;
 12'h2D4: rom_out <= 8'h00;
 12'h2D5: rom_out <= 8'h00;
 12'h2D6: rom_out <= 8'h00;
 12'h2D7: rom_out <= 8'h00;
 12'h2D8: rom_out <= 8'h00;
 12'h2D9: rom_out <= 8'h00;
 12'h2DA: rom_out <= 8'h00;
 12'h2DB: rom_out <= 8'h00;
 12'h2DC: rom_out <= 8'h00;
 12'h2DD: rom_out <= 8'h00;
 12'h2DE: rom_out <= 8'h00;
 12'h2DF: rom_out <= 8'h00;
 12'h2E0: rom_out <= 8'h00;
 12'h2E1: rom_out <= 8'h00;
 12'h2E2: rom_out <= 8'h00;
 12'h2E3: rom_out <= 8'h00;
 12'h2E4: rom_out <= 8'h00;
 12'h2E5: rom_out <= 8'h00;
 12'h2E6: rom_out <= 8'h00;
 12'h2E7: rom_out <= 8'h00;
 12'h2E8: rom_out <= 8'h00;
 12'h2E9: rom_out <= 8'h00;
 12'h2EA: rom_out <= 8'h00;
 12'h2EB: rom_out <= 8'h00;
 12'h2EC: rom_out <= 8'h00;
 12'h2ED: rom_out <= 8'h00;
 12'h2EE: rom_out <= 8'h00;
 12'h2EF: rom_out <= 8'h00;
 12'h2F0: rom_out <= 8'h00;
 12'h2F1: rom_out <= 8'h00;
 12'h2F2: rom_out <= 8'h00;
 12'h2F3: rom_out <= 8'h00;
 12'h2F4: rom_out <= 8'h00;
 12'h2F5: rom_out <= 8'h00;
 12'h2F6: rom_out <= 8'h00;
 12'h2F7: rom_out <= 8'h00;
 12'h2F8: rom_out <= 8'h00;
 12'h2F9: rom_out <= 8'h00;
 12'h2FA: rom_out <= 8'h00;
 12'h2FB: rom_out <= 8'h00;
 12'h2FC: rom_out <= 8'h00;
 12'h2FD: rom_out <= 8'h00;
 12'h2FE: rom_out <= 8'h00;
 12'h2FF: rom_out <= 8'h00;
  default: rom_out <= 8'h00;
	
	endcase
end

endmodule