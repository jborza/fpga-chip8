module dummy_rom(
	input wire [11:0] read_address,
	output reg [7:0] rom_out
);

always @* begin
	case (read_address)
		 'h200: rom_out <= 8'h00;
 'h201: rom_out <= 8'hE0;
 'h202: rom_out <= 8'hA2;
 'h203: rom_out <= 8'h2A;
 'h204: rom_out <= 8'h60;
 'h205: rom_out <= 8'h0C;
 'h206: rom_out <= 8'h61;
 'h207: rom_out <= 8'h08;
 'h208: rom_out <= 8'hD0;
 'h209: rom_out <= 8'h1F;
 'h20A: rom_out <= 8'h70;
 'h20B: rom_out <= 8'h09;
 'h20C: rom_out <= 8'hA2;
 'h20D: rom_out <= 8'h39;
 'h20E: rom_out <= 8'hD0;
 'h20F: rom_out <= 8'h1F;
 'h210: rom_out <= 8'hA2;
 'h211: rom_out <= 8'h48;
 'h212: rom_out <= 8'h70;
 'h213: rom_out <= 8'h08;
 'h214: rom_out <= 8'hD0;
 'h215: rom_out <= 8'h1F;
 'h216: rom_out <= 8'h70;
 'h217: rom_out <= 8'h04;
 'h218: rom_out <= 8'hA2;
 'h219: rom_out <= 8'h57;
 'h21A: rom_out <= 8'hD0;
 'h21B: rom_out <= 8'h1F;
 'h21C: rom_out <= 8'h70;
 'h21D: rom_out <= 8'h08;
 'h21E: rom_out <= 8'hA2;
 'h21F: rom_out <= 8'h66;
 'h220: rom_out <= 8'hD0;
 'h221: rom_out <= 8'h1F;
 'h222: rom_out <= 8'h70;
 'h223: rom_out <= 8'h08;
 'h224: rom_out <= 8'hA2;
 'h225: rom_out <= 8'h75;
 'h226: rom_out <= 8'hD0;
 'h227: rom_out <= 8'h1F;
 'h228: rom_out <= 8'h12;
 'h229: rom_out <= 8'h28;
 'h22A: rom_out <= 8'hFF;
 'h22B: rom_out <= 8'h00;
 'h22C: rom_out <= 8'hFF;
 'h22D: rom_out <= 8'h00;
 'h22E: rom_out <= 8'h3C;
 'h22F: rom_out <= 8'h00;
 'h230: rom_out <= 8'h3C;
 'h231: rom_out <= 8'h00;
 'h232: rom_out <= 8'h3C;
 'h233: rom_out <= 8'h00;
 'h234: rom_out <= 8'h3C;
 'h235: rom_out <= 8'h00;
 'h236: rom_out <= 8'hFF;
 'h237: rom_out <= 8'h00;
 'h238: rom_out <= 8'hFF;
 'h239: rom_out <= 8'hFF;
 'h23A: rom_out <= 8'h00;
 'h23B: rom_out <= 8'hFF;
 'h23C: rom_out <= 8'h00;
 'h23D: rom_out <= 8'h38;
 'h23E: rom_out <= 8'h00;
 'h23F: rom_out <= 8'h3F;
 'h240: rom_out <= 8'h00;
 'h241: rom_out <= 8'h3F;
 'h242: rom_out <= 8'h00;
 'h243: rom_out <= 8'h38;
 'h244: rom_out <= 8'h00;
 'h245: rom_out <= 8'hFF;
 'h246: rom_out <= 8'h00;
 'h247: rom_out <= 8'hFF;
 'h248: rom_out <= 8'h80;
 'h249: rom_out <= 8'h00;
 'h24A: rom_out <= 8'hE0;
 'h24B: rom_out <= 8'h00;
 'h24C: rom_out <= 8'hE0;
 'h24D: rom_out <= 8'h00;
 'h24E: rom_out <= 8'h80;
 'h24F: rom_out <= 8'h00;
 'h250: rom_out <= 8'h80;
 'h251: rom_out <= 8'h00;
 'h252: rom_out <= 8'hE0;
 'h253: rom_out <= 8'h00;
 'h254: rom_out <= 8'hE0;
 'h255: rom_out <= 8'h00;
 'h256: rom_out <= 8'h80;
 'h257: rom_out <= 8'hF8;
 'h258: rom_out <= 8'h00;
 'h259: rom_out <= 8'hFC;
 'h25A: rom_out <= 8'h00;
 'h25B: rom_out <= 8'h3E;
 'h25C: rom_out <= 8'h00;
 'h25D: rom_out <= 8'h3F;
 'h25E: rom_out <= 8'h00;
 'h25F: rom_out <= 8'h3B;
 'h260: rom_out <= 8'h00;
 'h261: rom_out <= 8'h39;
 'h262: rom_out <= 8'h00;
 'h263: rom_out <= 8'hF8;
 'h264: rom_out <= 8'h00;
 'h265: rom_out <= 8'hF8;
 'h266: rom_out <= 8'h03;
 'h267: rom_out <= 8'h00;
 'h268: rom_out <= 8'h07;
 'h269: rom_out <= 8'h00;
 'h26A: rom_out <= 8'h0F;
 'h26B: rom_out <= 8'h00;
 'h26C: rom_out <= 8'hBF;
 'h26D: rom_out <= 8'h00;
 'h26E: rom_out <= 8'hFB;
 'h26F: rom_out <= 8'h00;
 'h270: rom_out <= 8'hF3;
 'h271: rom_out <= 8'h00;
 'h272: rom_out <= 8'hE3;
 'h273: rom_out <= 8'h00;
 'h274: rom_out <= 8'h43;
 'h275: rom_out <= 8'hE0;
 'h276: rom_out <= 8'h00;
 'h277: rom_out <= 8'hE0;
 'h278: rom_out <= 8'h00;
 'h279: rom_out <= 8'h80;
 'h27A: rom_out <= 8'h00;
 'h27B: rom_out <= 8'h80;
 'h27C: rom_out <= 8'h00;
 'h27D: rom_out <= 8'h80;
 'h27E: rom_out <= 8'h00;
 'h27F: rom_out <= 8'h80;
 'h280: rom_out <= 8'h00;
 'h281: rom_out <= 8'hE0;
 'h282: rom_out <= 8'h00;
 'h283: rom_out <= 8'hE0;
 'h284: rom_out <= 8'h00;
 'h285: rom_out <= 8'h00;
 'h286: rom_out <= 8'h00;
 'h287: rom_out <= 8'h00;
 'h288: rom_out <= 8'h00;
 'h289: rom_out <= 8'h00;
 'h28A: rom_out <= 8'h00;
 'h28B: rom_out <= 8'h00;
 'h28C: rom_out <= 8'h00;
 'h28D: rom_out <= 8'h00;
 'h28E: rom_out <= 8'h00;
 'h28F: rom_out <= 8'h00;
 'h290: rom_out <= 8'h00;
 'h291: rom_out <= 8'h00;
 'h292: rom_out <= 8'h00;
 'h293: rom_out <= 8'h00;
 'h294: rom_out <= 8'h00;
 'h295: rom_out <= 8'h00;
 'h296: rom_out <= 8'h00;
 'h297: rom_out <= 8'h00;
 'h298: rom_out <= 8'h00;
 'h299: rom_out <= 8'h00;
 'h29A: rom_out <= 8'h00;
 'h29B: rom_out <= 8'h00;
 'h29C: rom_out <= 8'h00;
 'h29D: rom_out <= 8'h00;
 'h29E: rom_out <= 8'h00;
 'h29F: rom_out <= 8'h00;
 'h2A0: rom_out <= 8'h00;
 'h2A1: rom_out <= 8'h00;
 'h2A2: rom_out <= 8'h00;
 'h2A3: rom_out <= 8'h00;
 'h2A4: rom_out <= 8'h00;
 'h2A5: rom_out <= 8'h00;
 'h2A6: rom_out <= 8'h00;
 'h2A7: rom_out <= 8'h00;
 'h2A8: rom_out <= 8'h00;
 'h2A9: rom_out <= 8'h00;
 'h2AA: rom_out <= 8'h00;
 'h2AB: rom_out <= 8'h00;
 'h2AC: rom_out <= 8'h00;
 'h2AD: rom_out <= 8'h00;
 'h2AE: rom_out <= 8'h00;
 'h2AF: rom_out <= 8'h00;
 'h2B0: rom_out <= 8'h00;
 'h2B1: rom_out <= 8'h00;
 'h2B2: rom_out <= 8'h00;
 'h2B3: rom_out <= 8'h00;
 'h2B4: rom_out <= 8'h00;
 'h2B5: rom_out <= 8'h00;
 'h2B6: rom_out <= 8'h00;
 'h2B7: rom_out <= 8'h00;
 'h2B8: rom_out <= 8'h00;
 'h2B9: rom_out <= 8'h00;
 'h2BA: rom_out <= 8'h00;
 'h2BB: rom_out <= 8'h00;
 'h2BC: rom_out <= 8'h00;
 'h2BD: rom_out <= 8'h00;
 'h2BE: rom_out <= 8'h00;
 'h2BF: rom_out <= 8'h00;
 'h2C0: rom_out <= 8'h00;
 'h2C1: rom_out <= 8'h00;
 'h2C2: rom_out <= 8'h00;
 'h2C3: rom_out <= 8'h00;
 'h2C4: rom_out <= 8'h00;
 'h2C5: rom_out <= 8'h00;
 'h2C6: rom_out <= 8'h00;
 'h2C7: rom_out <= 8'h00;
 'h2C8: rom_out <= 8'h00;
 'h2C9: rom_out <= 8'h00;
 'h2CA: rom_out <= 8'h00;
 'h2CB: rom_out <= 8'h00;
 'h2CC: rom_out <= 8'h00;
 'h2CD: rom_out <= 8'h00;
 'h2CE: rom_out <= 8'h00;
 'h2CF: rom_out <= 8'h00;
 'h2D0: rom_out <= 8'h00;
 'h2D1: rom_out <= 8'h00;
 'h2D2: rom_out <= 8'h00;
 'h2D3: rom_out <= 8'h00;
 'h2D4: rom_out <= 8'h00;
 'h2D5: rom_out <= 8'h00;
 'h2D6: rom_out <= 8'h00;
 'h2D7: rom_out <= 8'h00;
 'h2D8: rom_out <= 8'h00;
 'h2D9: rom_out <= 8'h00;
 'h2DA: rom_out <= 8'h00;
 'h2DB: rom_out <= 8'h00;
 'h2DC: rom_out <= 8'h00;
 'h2DD: rom_out <= 8'h00;
 'h2DE: rom_out <= 8'h00;
 'h2DF: rom_out <= 8'h00;
 'h2E0: rom_out <= 8'h00;
 'h2E1: rom_out <= 8'h00;
 'h2E2: rom_out <= 8'h00;
 'h2E3: rom_out <= 8'h00;
 'h2E4: rom_out <= 8'h00;
 'h2E5: rom_out <= 8'h00;
 'h2E6: rom_out <= 8'h00;
 'h2E7: rom_out <= 8'h00;
 'h2E8: rom_out <= 8'h00;
 'h2E9: rom_out <= 8'h00;
 'h2EA: rom_out <= 8'h00;
 'h2EB: rom_out <= 8'h00;
 'h2EC: rom_out <= 8'h00;
 'h2ED: rom_out <= 8'h00;
 'h2EE: rom_out <= 8'h00;
 'h2EF: rom_out <= 8'h00;
 'h2F0: rom_out <= 8'h00;
 'h2F1: rom_out <= 8'h00;
 'h2F2: rom_out <= 8'h00;
 'h2F3: rom_out <= 8'h00;
 'h2F4: rom_out <= 8'h00;
 'h2F5: rom_out <= 8'h00;
 'h2F6: rom_out <= 8'h00;
 'h2F7: rom_out <= 8'h00;
 'h2F8: rom_out <= 8'h00;
 'h2F9: rom_out <= 8'h00;
 'h2FA: rom_out <= 8'h00;
 'h2FB: rom_out <= 8'h00;
 'h2FC: rom_out <= 8'h00;
 'h2FD: rom_out <= 8'h00;
 'h2FE: rom_out <= 8'h00;
 'h2FF: rom_out <= 8'h00;
  default: rom_out <= 8'h00;
	
	endcase
end

endmodule